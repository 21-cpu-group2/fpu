`default_nettype none
module fsqrt (
    input wire [31:0] op,
    output reg [31:0] result,
    input wire clk,
    input wire reset,
    output reg ready
);

reg [35:0] ram_read;
wire [23:0] ram_main;
wire [12:0] ram_grad;
assign ram_main = {1'b1, ram_read[35:13]};
assign ram_grad = ram_read[12:0];

reg [35:0] ram [1023:0];

reg [7:0] exp2;
reg [13:0] res;

reg [7:0] exp3;
reg [26:0] grad_mul_res;
reg [23:0] frac;

always @(posedge clk) begin
    if (~reset) begin
        result <= 32'd0;
        ready <= 1'b0;
        exp2 <= 8'd0;
		exp3 <= 8'd0;
		grad_mul_res <= 27'd0;
		frac <= 24'd0;
		ram[0] <= 36'b011010100000100111100110101101001110;
		ram[1] <= 36'b011010100110010001011100101101001100;
		ram[2] <= 36'b011010101011111010111110101101001001;
		ram[3] <= 36'b011010110001100100001000101101000110;
		ram[4] <= 36'b011010110111001100111010101101000011;
		ram[5] <= 36'b011010111100110101011000101101000000;
		ram[6] <= 36'b011011000010011101100000101100111110;
		ram[7] <= 36'b011011001000000101010000101100111011;
		ram[8] <= 36'b011011001101101100101010101100111000;
		ram[9] <= 36'b011011010011010011110000101100110101;
		ram[10] <= 36'b011011011000111010011110101100110011;
		ram[11] <= 36'b011011011110100000110110101100110000;
		ram[12] <= 36'b011011100100000110111000101100101101;
		ram[13] <= 36'b011011101001101100100110101100101010;
		ram[14] <= 36'b011011101111010001111100101100101000;
		ram[15] <= 36'b011011110100110110111110101100100101;
		ram[16] <= 36'b011011111010011011101010101100100010;
		ram[17] <= 36'b011100000000000000000000101100100000;
		ram[18] <= 36'b011100000101100100000000101100011101;
		ram[19] <= 36'b011100001011000111101010101100011010;
		ram[20] <= 36'b011100010000101011000000101100011000;
		ram[21] <= 36'b011100010110001110000000101100010101;
		ram[22] <= 36'b011100011011110000101010101100010010;
		ram[23] <= 36'b011100100001010011000000101100010000;
		ram[24] <= 36'b011100100110110101000000101100001101;
		ram[25] <= 36'b011100101100010110101100101100001010;
		ram[26] <= 36'b011100110001111000000010101100001000;
		ram[27] <= 36'b011100110111011001000100101100000101;
		ram[28] <= 36'b011100111100111001110000101100000010;
		ram[29] <= 36'b011101000010011010000110101100000000;
		ram[30] <= 36'b011101000111111010001010101011111101;
		ram[31] <= 36'b011101001101011001110110101011111011;
		ram[32] <= 36'b011101010010111001010000101011111000;
		ram[33] <= 36'b011101011000011000010100101011110101;
		ram[34] <= 36'b011101011101110111000100101011110011;
		ram[35] <= 36'b011101100011010101100000101011110000;
		ram[36] <= 36'b011101101000110011100110101011101110;
		ram[37] <= 36'b011101101110010001011000101011101011;
		ram[38] <= 36'b011101110011101110110110101011101001;
		ram[39] <= 36'b011101111001001100000000101011100110;
		ram[40] <= 36'b011101111110101000110100101011100100;
		ram[41] <= 36'b011110000100000101010110101011100001;
		ram[42] <= 36'b011110001001100001100010101011011111;
		ram[43] <= 36'b011110001110111101011100101011011100;
		ram[44] <= 36'b011110010100011001000000101011011010;
		ram[45] <= 36'b011110011001110100010010101011010111;
		ram[46] <= 36'b011110011111001111001110101011010101;
		ram[47] <= 36'b011110100100101001110110101011010010;
		ram[48] <= 36'b011110101010000100001100101011010000;
		ram[49] <= 36'b011110101111011110001110101011001101;
		ram[50] <= 36'b011110110100110111111100101011001011;
		ram[51] <= 36'b011110111010010001010100101011001000;
		ram[52] <= 36'b011110111111101010011100101011000110;
		ram[53] <= 36'b011111000101000011001110101011000011;
		ram[54] <= 36'b011111001010011011101110101011000001;
		ram[55] <= 36'b011111001111110011111000101010111111;
		ram[56] <= 36'b011111010101001011110010101010111100;
		ram[57] <= 36'b011111011010100011010110101010111010;
		ram[58] <= 36'b011111011111111010101000101010110111;
		ram[59] <= 36'b011111100101010001100110101010110101;
		ram[60] <= 36'b011111101010101000010010101010110011;
		ram[61] <= 36'b011111101111111110101010101010110000;
		ram[62] <= 36'b011111110101010100101110101010101110;
		ram[63] <= 36'b011111111010101010100000101010101011;
		ram[64] <= 36'b100000000000000000000000101010101001;
		ram[65] <= 36'b100000000101010101001010101010100111;
		ram[66] <= 36'b100000001010101010000100101010100100;
		ram[67] <= 36'b100000001111111110101010101010100010;
		ram[68] <= 36'b100000010101010010111110101010100000;
		ram[69] <= 36'b100000011010100110111110101010011101;
		ram[70] <= 36'b100000011111111010101100101010011011;
		ram[71] <= 36'b100000100101001110000110101010011001;
		ram[72] <= 36'b100000101010100001010000101010010110;
		ram[73] <= 36'b100000101111110100000100101010010100;
		ram[74] <= 36'b100000110101000110101000101010010010;
		ram[75] <= 36'b100000111010011000111010101010001111;
		ram[76] <= 36'b100000111111101010111000101010001101;
		ram[77] <= 36'b100001000100111100100100101010001011;
		ram[78] <= 36'b100001001010001101111110101010001000;
		ram[79] <= 36'b100001001111011111000110101010000110;
		ram[80] <= 36'b100001010100101111111010101010000100;
		ram[81] <= 36'b100001011010000000011110101010000010;
		ram[82] <= 36'b100001011111010000101110101001111111;
		ram[83] <= 36'b100001100100100000101100101001111101;
		ram[84] <= 36'b100001101001110000011010101001111011;
		ram[85] <= 36'b100001101110111111110100101001111001;
		ram[86] <= 36'b100001110100001110111100101001110110;
		ram[87] <= 36'b100001111001011101110100101001110100;
		ram[88] <= 36'b100001111110101100011000101001110010;
		ram[89] <= 36'b100010000011111010101100101001110000;
		ram[90] <= 36'b100010001001001000101100101001101101;
		ram[91] <= 36'b100010001110010110011100101001101011;
		ram[92] <= 36'b100010010011100011111010101001101001;
		ram[93] <= 36'b100010011000110001000110101001100111;
		ram[94] <= 36'b100010011101111110000000101001100101;
		ram[95] <= 36'b100010100011001010101010101001100010;
		ram[96] <= 36'b100010101000010111000010101001100000;
		ram[97] <= 36'b100010101101100011001000101001011110;
		ram[98] <= 36'b100010110010101110111100101001011100;
		ram[99] <= 36'b100010110111111010011110101001011010;
		ram[100] <= 36'b100010111101000101110000101001011000;
		ram[101] <= 36'b100011000010010000110010101001010101;
		ram[102] <= 36'b100011000111011011100000101001010011;
		ram[103] <= 36'b100011001100100101111110101001010001;
		ram[104] <= 36'b100011010001110000001010101001001111;
		ram[105] <= 36'b100011010110111010000110101001001101;
		ram[106] <= 36'b100011011100000011110010101001001011;
		ram[107] <= 36'b100011100001001101001010101001001001;
		ram[108] <= 36'b100011100110010110010010101001000110;
		ram[109] <= 36'b100011101011011111001010101001000100;
		ram[110] <= 36'b100011110000100111110000101001000010;
		ram[111] <= 36'b100011110101110000000110101001000000;
		ram[112] <= 36'b100011111010111000001100101000111110;
		ram[113] <= 36'b100100000000000000000000101000111100;
		ram[114] <= 36'b100100000101000111100010101000111010;
		ram[115] <= 36'b100100001010001110110100101000111000;
		ram[116] <= 36'b100100001111010101110110101000110110;
		ram[117] <= 36'b100100010100011100101000101000110100;
		ram[118] <= 36'b100100011001100011001000101000110001;
		ram[119] <= 36'b100100011110101001011000101000101111;
		ram[120] <= 36'b100100100011101111010110101000101101;
		ram[121] <= 36'b100100101000110101000110101000101011;
		ram[122] <= 36'b100100101101111010100100101000101001;
		ram[123] <= 36'b100100110010111111110010101000100111;
		ram[124] <= 36'b100100111000000100110000101000100101;
		ram[125] <= 36'b100100111101001001011100101000100011;
		ram[126] <= 36'b100101000010001101111010101000100001;
		ram[127] <= 36'b100101000111010010000110101000011111;
		ram[128] <= 36'b100101001100010110000010101000011101;
		ram[129] <= 36'b100101010001011001101110101000011011;
		ram[130] <= 36'b100101010110011101001010101000011001;
		ram[131] <= 36'b100101011011100000010110101000010111;
		ram[132] <= 36'b100101100000100011010010101000010101;
		ram[133] <= 36'b100101100101100101111110101000010011;
		ram[134] <= 36'b100101101010101000011010101000010001;
		ram[135] <= 36'b100101101111101010100110101000001111;
		ram[136] <= 36'b100101110100101100100010101000001101;
		ram[137] <= 36'b100101111001101110001110101000001011;
		ram[138] <= 36'b100101111110101111101010101000001001;
		ram[139] <= 36'b100110000011110000110110101000000111;
		ram[140] <= 36'b100110001000110001110100101000000101;
		ram[141] <= 36'b100110001101110010100000101000000011;
		ram[142] <= 36'b100110010010110010111110101000000001;
		ram[143] <= 36'b100110010111110011001010100111111111;
		ram[144] <= 36'b100110011100110011001000100111111101;
		ram[145] <= 36'b100110100001110010110110100111111011;
		ram[146] <= 36'b100110100110110010010110100111111001;
		ram[147] <= 36'b100110101011110001100100100111110111;
		ram[148] <= 36'b100110110000110000100100100111110110;
		ram[149] <= 36'b100110110101101111010100100111110100;
		ram[150] <= 36'b100110111010101101110110100111110010;
		ram[151] <= 36'b100110111111101100000110100111110000;
		ram[152] <= 36'b100111000100101010001000100111101110;
		ram[153] <= 36'b100111001001100111111100100111101100;
		ram[154] <= 36'b100111001110100101011110100111101010;
		ram[155] <= 36'b100111010011100010110010100111101000;
		ram[156] <= 36'b100111011000011111111000100111100110;
		ram[157] <= 36'b100111011101011100101110100111100100;
		ram[158] <= 36'b100111100010011001010100100111100010;
		ram[159] <= 36'b100111100111010101101100100111100001;
		ram[160] <= 36'b100111101100010001110100100111011111;
		ram[161] <= 36'b100111110001001101101100100111011101;
		ram[162] <= 36'b100111110110001001011000100111011011;
		ram[163] <= 36'b100111111011000100110010100111011001;
		ram[164] <= 36'b101000000000000000000000100111010111;
		ram[165] <= 36'b101000000100111010111100100111010101;
		ram[166] <= 36'b101000001001110101101100100111010011;
		ram[167] <= 36'b101000001110110000001010100111010010;
		ram[168] <= 36'b101000010011101010011100100111010000;
		ram[169] <= 36'b101000011000100100011110100111001110;
		ram[170] <= 36'b101000011101011110010010100111001100;
		ram[171] <= 36'b101000100010010111110110100111001010;
		ram[172] <= 36'b101000100111010001001100100111001000;
		ram[173] <= 36'b101000101100001010010100100111000111;
		ram[174] <= 36'b101000110001000011001100100111000101;
		ram[175] <= 36'b101000110101111011110110100111000011;
		ram[176] <= 36'b101000111010110100010010100111000001;
		ram[177] <= 36'b101000111111101100011110100110111111;
		ram[178] <= 36'b101001000100100100011110100110111110;
		ram[179] <= 36'b101001001001011100001110100110111100;
		ram[180] <= 36'b101001001110010011101110100110111010;
		ram[181] <= 36'b101001010011001011000010100110111000;
		ram[182] <= 36'b101001011000000010001000100110110110;
		ram[183] <= 36'b101001011100111000111110100110110101;
		ram[184] <= 36'b101001100001101111100110100110110011;
		ram[185] <= 36'b101001100110100110000000100110110001;
		ram[186] <= 36'b101001101011011100001100100110101111;
		ram[187] <= 36'b101001110000010010001000100110101101;
		ram[188] <= 36'b101001110101000111111000100110101100;
		ram[189] <= 36'b101001111001111101011010100110101010;
		ram[190] <= 36'b101001111110110010101100100110101000;
		ram[191] <= 36'b101010000011100111110010100110100110;
		ram[192] <= 36'b101010001000011100101000100110100101;
		ram[193] <= 36'b101010001101010001010010100110100011;
		ram[194] <= 36'b101010010010000101101100100110100001;
		ram[195] <= 36'b101010010110111001111000100110011111;
		ram[196] <= 36'b101010011011101101111000100110011110;
		ram[197] <= 36'b101010100000100001101000100110011100;
		ram[198] <= 36'b101010100101010101001100100110011010;
		ram[199] <= 36'b101010101010001000100010100110011000;
		ram[200] <= 36'b101010101110111011101000100110010111;
		ram[201] <= 36'b101010110011101110100010100110010101;
		ram[202] <= 36'b101010111000100001001110100110010011;
		ram[203] <= 36'b101010111101010011101100100110010010;
		ram[204] <= 36'b101011000010000101111100100110010000;
		ram[205] <= 36'b101011000110111000000000100110001110;
		ram[206] <= 36'b101011001011101001110100100110001100;
		ram[207] <= 36'b101011010000011011011100100110001011;
		ram[208] <= 36'b101011010101001100110110100110001001;
		ram[209] <= 36'b101011011001111110000010100110000111;
		ram[210] <= 36'b101011011110101111000000100110000110;
		ram[211] <= 36'b101011100011011111110010100110000100;
		ram[212] <= 36'b101011101000010000010110100110000010;
		ram[213] <= 36'b101011101101000000101100100110000001;
		ram[214] <= 36'b101011110001110000110100100101111111;
		ram[215] <= 36'b101011110110100000110000100101111101;
		ram[216] <= 36'b101011111011010000011110100101111100;
		ram[217] <= 36'b101100000000000000000000100101111010;
		ram[218] <= 36'b101100000100101111010010100101111000;
		ram[219] <= 36'b101100001001011110011000100101110111;
		ram[220] <= 36'b101100001110001101010010100101110101;
		ram[221] <= 36'b101100010010111011111110100101110011;
		ram[222] <= 36'b101100010111101010011100100101110010;
		ram[223] <= 36'b101100011100011000101100100101110000;
		ram[224] <= 36'b101100100001000110110000100101101110;
		ram[225] <= 36'b101100100101110100101000100101101101;
		ram[226] <= 36'b101100101010100010010010100101101011;
		ram[227] <= 36'b101100101111001111101110100101101001;
		ram[228] <= 36'b101100110011111100111110100101101000;
		ram[229] <= 36'b101100111000101010000000100101100110;
		ram[230] <= 36'b101100111101010110110110100101100101;
		ram[231] <= 36'b101101000010000011100000100101100011;
		ram[232] <= 36'b101101000110101111111100100101100001;
		ram[233] <= 36'b101101001011011100001010100101100000;
		ram[234] <= 36'b101101010000001000001100100101011110;
		ram[235] <= 36'b101101010100110100000010100101011101;
		ram[236] <= 36'b101101011001011111101010100101011011;
		ram[237] <= 36'b101101011110001011000100100101011001;
		ram[238] <= 36'b101101100010110110010100100101011000;
		ram[239] <= 36'b101101100111100001010110100101010110;
		ram[240] <= 36'b101101101100001100001010100101010101;
		ram[241] <= 36'b101101110000110110110010100101010011;
		ram[242] <= 36'b101101110101100001001110100101010001;
		ram[243] <= 36'b101101111010001011011110100101010000;
		ram[244] <= 36'b101101111110110101100000100101001110;
		ram[245] <= 36'b101110000011011111010110100101001101;
		ram[246] <= 36'b101110001000001001000000100101001011;
		ram[247] <= 36'b101110001100110010011100100101001010;
		ram[248] <= 36'b101110010001011011101100100101001000;
		ram[249] <= 36'b101110010110000100110000100101000110;
		ram[250] <= 36'b101110011010101101101000100101000101;
		ram[251] <= 36'b101110011111010110010010100101000011;
		ram[252] <= 36'b101110100011111110110000100101000010;
		ram[253] <= 36'b101110101000100111000010100101000000;
		ram[254] <= 36'b101110101101001111001000100100111111;
		ram[255] <= 36'b101110110001110111000000100100111101;
		ram[256] <= 36'b101110110110011110101110100100111100;
		ram[257] <= 36'b101110111011000110001110100100111010;
		ram[258] <= 36'b101110111111101101100010100100111000;
		ram[259] <= 36'b101111000100010100101010100100110111;
		ram[260] <= 36'b101111001000111011100110100100110101;
		ram[261] <= 36'b101111001101100010010110100100110100;
		ram[262] <= 36'b101111010010001000111000100100110010;
		ram[263] <= 36'b101111010110101111010000100100110001;
		ram[264] <= 36'b101111011011010101011010100100101111;
		ram[265] <= 36'b101111011111111011011010100100101110;
		ram[266] <= 36'b101111100100100001001100100100101100;
		ram[267] <= 36'b101111101001000110110010100100101011;
		ram[268] <= 36'b101111101101101100001100100100101001;
		ram[269] <= 36'b101111110010010001011100100100101000;
		ram[270] <= 36'b101111110110110110011110100100100110;
		ram[271] <= 36'b101111111011011011010100100100100101;
		ram[272] <= 36'b110000000000000000000000100100100011;
		ram[273] <= 36'b110000000100100100011110100100100010;
		ram[274] <= 36'b110000001001001000110000100100100000;
		ram[275] <= 36'b110000001101101100111000100100011111;
		ram[276] <= 36'b110000010010010000110010100100011101;
		ram[277] <= 36'b110000010110110100100010100100011100;
		ram[278] <= 36'b110000011011011000000100100100011010;
		ram[279] <= 36'b110000011111111011011100100100011001;
		ram[280] <= 36'b110000100100011110101000100100010111;
		ram[281] <= 36'b110000101001000001101000100100010110;
		ram[282] <= 36'b110000101101100100011100100100010101;
		ram[283] <= 36'b110000110010000111000100100100010011;
		ram[284] <= 36'b110000110110101001100000100100010010;
		ram[285] <= 36'b110000111011001011110010100100010000;
		ram[286] <= 36'b110000111111101101111000100100001111;
		ram[287] <= 36'b110001000100001111110000100100001101;
		ram[288] <= 36'b110001001000110001100000100100001100;
		ram[289] <= 36'b110001001101010011000010100100001010;
		ram[290] <= 36'b110001010001110100011000100100001001;
		ram[291] <= 36'b110001010110010101100100100100000111;
		ram[292] <= 36'b110001011010110110100100100100000110;
		ram[293] <= 36'b110001011111010111011000100100000101;
		ram[294] <= 36'b110001100011111000000010100100000011;
		ram[295] <= 36'b110001101000011000100000100100000010;
		ram[296] <= 36'b110001101100111000110010100100000000;
		ram[297] <= 36'b110001110001011000111000100011111111;
		ram[298] <= 36'b110001110101111000110100100011111101;
		ram[299] <= 36'b110001111010011000100100100011111100;
		ram[300] <= 36'b110001111110111000001000100011111011;
		ram[301] <= 36'b110010000011010111100000100011111001;
		ram[302] <= 36'b110010000111110110101110100011111000;
		ram[303] <= 36'b110010001100010101110010100011110110;
		ram[304] <= 36'b110010010000110100101000100011110101;
		ram[305] <= 36'b110010010101010011010100100011110100;
		ram[306] <= 36'b110010011001110001110110100011110010;
		ram[307] <= 36'b110010011110010000001100100011110001;
		ram[308] <= 36'b110010100010101110010110100011101111;
		ram[309] <= 36'b110010100111001100010110100011101110;
		ram[310] <= 36'b110010101011101010001010100011101101;
		ram[311] <= 36'b110010110000000111110010100011101011;
		ram[312] <= 36'b110010110100100101010000100011101010;
		ram[313] <= 36'b110010111001000010100100100011101000;
		ram[314] <= 36'b110010111101011111101100100011100111;
		ram[315] <= 36'b110011000001111100101000100011100110;
		ram[316] <= 36'b110011000110011001011010100011100100;
		ram[317] <= 36'b110011001010110110000000100011100011;
		ram[318] <= 36'b110011001111010010011100100011100010;
		ram[319] <= 36'b110011010011101110101110100011100000;
		ram[320] <= 36'b110011011000001010110100100011011111;
		ram[321] <= 36'b110011011100100110101110100011011110;
		ram[322] <= 36'b110011100001000010011110100011011100;
		ram[323] <= 36'b110011100101011110000100100011011011;
		ram[324] <= 36'b110011101001111001011110100011011001;
		ram[325] <= 36'b110011101110010100101110100011011000;
		ram[326] <= 36'b110011110010101111110010100011010111;
		ram[327] <= 36'b110011110111001010101100100011010101;
		ram[328] <= 36'b110011111011100101011010100011010100;
		ram[329] <= 36'b110100000000000000000000100011010011;
		ram[330] <= 36'b110100000100011010011000100011010001;
		ram[331] <= 36'b110100001000110100101000100011010000;
		ram[332] <= 36'b110100001101001110101100100011001111;
		ram[333] <= 36'b110100010001101000100100100011001101;
		ram[334] <= 36'b110100010110000010010100100011001100;
		ram[335] <= 36'b110100011010011011111000100011001011;
		ram[336] <= 36'b110100011110110101010010100011001001;
		ram[337] <= 36'b110100100011001110100000100011001000;
		ram[338] <= 36'b110100100111100111100100100011000111;
		ram[339] <= 36'b110100101100000000011110100011000101;
		ram[340] <= 36'b110100110000011001001100100011000100;
		ram[341] <= 36'b110100110100110001110010100011000011;
		ram[342] <= 36'b110100111001001010001100100011000001;
		ram[343] <= 36'b110100111101100010011010100011000000;
		ram[344] <= 36'b110101000001111010100000100010111111;
		ram[345] <= 36'b110101000110010010011010100010111110;
		ram[346] <= 36'b110101001010101010001010100010111100;
		ram[347] <= 36'b110101001111000001110000100010111011;
		ram[348] <= 36'b110101010011011001001100100010111010;
		ram[349] <= 36'b110101010111110000011100100010111000;
		ram[350] <= 36'b110101011100000111100010100010110111;
		ram[351] <= 36'b110101100000011110100000100010110110;
		ram[352] <= 36'b110101100100110101010000100010110100;
		ram[353] <= 36'b110101101001001011111000100010110011;
		ram[354] <= 36'b110101101101100010010110100010110010;
		ram[355] <= 36'b110101110001111000101000100010110001;
		ram[356] <= 36'b110101110110001110110010100010101111;
		ram[357] <= 36'b110101111010100100110000100010101110;
		ram[358] <= 36'b110101111110111010100100100010101101;
		ram[359] <= 36'b110110000011010000001110100010101011;
		ram[360] <= 36'b110110000111100101101110100010101010;
		ram[361] <= 36'b110110001011111011000010100010101001;
		ram[362] <= 36'b110110010000010000001110100010101000;
		ram[363] <= 36'b110110010100100101010000100010100110;
		ram[364] <= 36'b110110011000111010000110100010100101;
		ram[365] <= 36'b110110011101001110110100100010100100;
		ram[366] <= 36'b110110100001100011010110100010100011;
		ram[367] <= 36'b110110100101110111110000100010100001;
		ram[368] <= 36'b110110101010001011111110100010100000;
		ram[369] <= 36'b110110101110100000000010100010011111;
		ram[370] <= 36'b110110110010110011111110100010011110;
		ram[371] <= 36'b110110110111000111101110100010011100;
		ram[372] <= 36'b110110111011011011010100100010011011;
		ram[373] <= 36'b110110111111101110110010100010011010;
		ram[374] <= 36'b110111000100000010000100100010011001;
		ram[375] <= 36'b110111001000010101001110100010010111;
		ram[376] <= 36'b110111001100101000001100100010010110;
		ram[377] <= 36'b110111010000111011000010100010010101;
		ram[378] <= 36'b110111010101001101101100100010010100;
		ram[379] <= 36'b110111011001100000001110100010010010;
		ram[380] <= 36'b110111011101110010100100100010010001;
		ram[381] <= 36'b110111100010000100110010100010010000;
		ram[382] <= 36'b110111100110010110110110100010001111;
		ram[383] <= 36'b110111101010101000110000100010001110;
		ram[384] <= 36'b110111101110111010100000100010001100;
		ram[385] <= 36'b110111110011001100000110100010001011;
		ram[386] <= 36'b110111110111011101100100100010001010;
		ram[387] <= 36'b110111111011101110110110100010001001;
		ram[388] <= 36'b111000000000000000000000100010000111;
		ram[389] <= 36'b111000000100010000111110100010000110;
		ram[390] <= 36'b111000001000100001110100100010000101;
		ram[391] <= 36'b111000001100110010100000100010000100;
		ram[392] <= 36'b111000010001000011000010100010000011;
		ram[393] <= 36'b111000010101010011011100100010000001;
		ram[394] <= 36'b111000011001100011101010100010000000;
		ram[395] <= 36'b111000011101110011110000100001111111;
		ram[396] <= 36'b111000100010000011101100100001111110;
		ram[397] <= 36'b111000100110010011011110100001111101;
		ram[398] <= 36'b111000101010100011000110100001111011;
		ram[399] <= 36'b111000101110110010100110100001111010;
		ram[400] <= 36'b111000110011000001111100100001111001;
		ram[401] <= 36'b111000110111010001001000100001111000;
		ram[402] <= 36'b111000111011100000001010100001110111;
		ram[403] <= 36'b111000111111101111000100100001110101;
		ram[404] <= 36'b111001000011111101110100100001110100;
		ram[405] <= 36'b111001001000001100011010100001110011;
		ram[406] <= 36'b111001001100011010110110100001110010;
		ram[407] <= 36'b111001010000101001001010100001110001;
		ram[408] <= 36'b111001010100110111010100100001110000;
		ram[409] <= 36'b111001011001000101010100100001101110;
		ram[410] <= 36'b111001011101010011001100100001101101;
		ram[411] <= 36'b111001100001100000111010100001101100;
		ram[412] <= 36'b111001100101101110011110100001101011;
		ram[413] <= 36'b111001101001111011111010100001101010;
		ram[414] <= 36'b111001101110001001001010100001101001;
		ram[415] <= 36'b111001110010010110010100100001100111;
		ram[416] <= 36'b111001110110100011010010100001100110;
		ram[417] <= 36'b111001111010110000001000100001100101;
		ram[418] <= 36'b111001111110111100110110100001100100;
		ram[419] <= 36'b111010000011001001011000100001100011;
		ram[420] <= 36'b111010000111010101110010100001100010;
		ram[421] <= 36'b111010001011100010000100100001100000;
		ram[422] <= 36'b111010001111101110001100100001011111;
		ram[423] <= 36'b111010010011111010001010100001011110;
		ram[424] <= 36'b111010011000000110000000100001011101;
		ram[425] <= 36'b111010011100010001101100100001011100;
		ram[426] <= 36'b111010100000011101010000100001011011;
		ram[427] <= 36'b111010100100101000101010100001011010;
		ram[428] <= 36'b111010101000110011111010100001011000;
		ram[429] <= 36'b111010101100111111000010100001010111;
		ram[430] <= 36'b111010110001001010000000100001010110;
		ram[431] <= 36'b111010110101010100110110100001010101;
		ram[432] <= 36'b111010111001011111100100100001010100;
		ram[433] <= 36'b111010111101101010000110100001010011;
		ram[434] <= 36'b111011000001110100100010100001010010;
		ram[435] <= 36'b111011000101111110110100100001010001;
		ram[436] <= 36'b111011001010001000111100100001001111;
		ram[437] <= 36'b111011001110010010111100100001001110;
		ram[438] <= 36'b111011010010011100110010100001001101;
		ram[439] <= 36'b111011010110100110100000100001001100;
		ram[440] <= 36'b111011011010110000000100100001001011;
		ram[441] <= 36'b111011011110111001100000100001001010;
		ram[442] <= 36'b111011100011000010110100100001001001;
		ram[443] <= 36'b111011100111001011111110100001001000;
		ram[444] <= 36'b111011101011010100111110100001000111;
		ram[445] <= 36'b111011101111011101110110100001000101;
		ram[446] <= 36'b111011110011100110100110100001000100;
		ram[447] <= 36'b111011110111101111001100100001000011;
		ram[448] <= 36'b111011111011110111101010100001000010;
		ram[449] <= 36'b111100000000000000000000100001000001;
		ram[450] <= 36'b111100000100001000001100100001000000;
		ram[451] <= 36'b111100001000010000001110100000111111;
		ram[452] <= 36'b111100001100011000001010100000111110;
		ram[453] <= 36'b111100010000011111111010100000111101;
		ram[454] <= 36'b111100010100100111100100100000111100;
		ram[455] <= 36'b111100011000101111000100100000111010;
		ram[456] <= 36'b111100011100110110011100100000111001;
		ram[457] <= 36'b111100100000111101101010100000111000;
		ram[458] <= 36'b111100100101000100110000100000110111;
		ram[459] <= 36'b111100101001001011101110100000110110;
		ram[460] <= 36'b111100101101010010100100100000110101;
		ram[461] <= 36'b111100110001011001010000100000110100;
		ram[462] <= 36'b111100110101011111110100100000110011;
		ram[463] <= 36'b111100111001100110001110100000110010;
		ram[464] <= 36'b111100111101101100100000100000110001;
		ram[465] <= 36'b111101000001110010101010100000110000;
		ram[466] <= 36'b111101000101111000101100100000101111;
		ram[467] <= 36'b111101001001111110100100100000101110;
		ram[468] <= 36'b111101001110000100010100100000101100;
		ram[469] <= 36'b111101010010001001111100100000101011;
		ram[470] <= 36'b111101010110001111011010100000101010;
		ram[471] <= 36'b111101011010010100110000100000101001;
		ram[472] <= 36'b111101011110011001111110100000101000;
		ram[473] <= 36'b111101100010011111000100100000100111;
		ram[474] <= 36'b111101100110100100000010100000100110;
		ram[475] <= 36'b111101101010101000110110100000100101;
		ram[476] <= 36'b111101101110101101100010100000100100;
		ram[477] <= 36'b111101110010110010000110100000100011;
		ram[478] <= 36'b111101110110110110100000100000100010;
		ram[479] <= 36'b111101111010111010110100100000100001;
		ram[480] <= 36'b111101111110111110111110100000100000;
		ram[481] <= 36'b111110000011000011000000100000011111;
		ram[482] <= 36'b111110000111000110111010100000011110;
		ram[483] <= 36'b111110001011001010101010100000011101;
		ram[484] <= 36'b111110001111001110010100100000011100;
		ram[485] <= 36'b111110010011010001110100100000011011;
		ram[486] <= 36'b111110010111010101001100100000011001;
		ram[487] <= 36'b111110011011011000011100100000011000;
		ram[488] <= 36'b111110011111011011100100100000010111;
		ram[489] <= 36'b111110100011011110100010100000010110;
		ram[490] <= 36'b111110100111100001011010100000010101;
		ram[491] <= 36'b111110101011100100001000100000010100;
		ram[492] <= 36'b111110101111100110110000100000010011;
		ram[493] <= 36'b111110110011101001001110100000010010;
		ram[494] <= 36'b111110110111101011100100100000010001;
		ram[495] <= 36'b111110111011101101110010100000010000;
		ram[496] <= 36'b111110111111101111110110100000001111;
		ram[497] <= 36'b111111000011110001110100100000001110;
		ram[498] <= 36'b111111000111110011101010100000001101;
		ram[499] <= 36'b111111001011110101010110100000001100;
		ram[500] <= 36'b111111001111110110111100100000001011;
		ram[501] <= 36'b111111010011111000011000100000001010;
		ram[502] <= 36'b111111010111111001101110100000001001;
		ram[503] <= 36'b111111011011111010111010100000001000;
		ram[504] <= 36'b111111011111111011111110100000000111;
		ram[505] <= 36'b111111100011111100111010100000000110;
		ram[506] <= 36'b111111100111111101101110100000000101;
		ram[507] <= 36'b111111101011111110011010100000000100;
		ram[508] <= 36'b111111101111111110111110100000000011;
		ram[509] <= 36'b111111110011111111011010100000000010;
		ram[510] <= 36'b111111110111111111101110100000000001;
		ram[511] <= 36'b111111111011111111111010100000000000;
		ram[512] <= 36'b000000000000000000000001000000000000;
		ram[513] <= 36'b000000000011111111111000111111111100;
		ram[514] <= 36'b000000000111111111100000111111111000;
		ram[515] <= 36'b000000001011111110111000111111110100;
		ram[516] <= 36'b000000001111111110000000111111110000;
		ram[517] <= 36'b000000010011111100111000111111101100;
		ram[518] <= 36'b000000010111111011100000111111101000;
		ram[519] <= 36'b000000011011111001111010111111100100;
		ram[520] <= 36'b000000011111111000000010111111100000;
		ram[521] <= 36'b000000100011110101111100111111011100;
		ram[522] <= 36'b000000100111110011100110111111011000;
		ram[523] <= 36'b000000101011110001000010111111010100;
		ram[524] <= 36'b000000101111101110001100111111010000;
		ram[525] <= 36'b000000110011101011001000111111001100;
		ram[526] <= 36'b000000110111100111110100111111001001;
		ram[527] <= 36'b000000111011100100010000111111000101;
		ram[528] <= 36'b000000111111100000011110111111000001;
		ram[529] <= 36'b000001000011011100011100111110111101;
		ram[530] <= 36'b000001000111011000001100111110111001;
		ram[531] <= 36'b000001001011010011101100111110110110;
		ram[532] <= 36'b000001001111001110111100111110110010;
		ram[533] <= 36'b000001010011001001111110111110101110;
		ram[534] <= 36'b000001010111000100110000111110101010;
		ram[535] <= 36'b000001011010111111010100111110100110;
		ram[536] <= 36'b000001011110111001101000111110100011;
		ram[537] <= 36'b000001100010110011101110111110011111;
		ram[538] <= 36'b000001100110101101100100111110011011;
		ram[539] <= 36'b000001101010100111001100111110011000;
		ram[540] <= 36'b000001101110100000100100111110010100;
		ram[541] <= 36'b000001110010011001110000111110010000;
		ram[542] <= 36'b000001110110010010101010111110001101;
		ram[543] <= 36'b000001111010001011011000111110001001;
		ram[544] <= 36'b000001111110000011110110111110000101;
		ram[545] <= 36'b000010000001111100000100111110000010;
		ram[546] <= 36'b000010000101110100000110111101111110;
		ram[547] <= 36'b000010001001101011111000111101111010;
		ram[548] <= 36'b000010001101100011011100111101110111;
		ram[549] <= 36'b000010010001011010110010111101110011;
		ram[550] <= 36'b000010010101010001111000111101101111;
		ram[551] <= 36'b000010011001001000110010111101101100;
		ram[552] <= 36'b000010011100111111011100111101101000;
		ram[553] <= 36'b000010100000110101111000111101100101;
		ram[554] <= 36'b000010100100101100000110111101100001;
		ram[555] <= 36'b000010101000100010000110111101011110;
		ram[556] <= 36'b000010101100010111110110111101011010;
		ram[557] <= 36'b000010110000001101011010111101010111;
		ram[558] <= 36'b000010110100000010110000111101010011;
		ram[559] <= 36'b000010110111110111110110111101010000;
		ram[560] <= 36'b000010111011101100110000111101001100;
		ram[561] <= 36'b000010111111100001011010111101001001;
		ram[562] <= 36'b000011000011010101111000111101000101;
		ram[563] <= 36'b000011000111001010001000111101000010;
		ram[564] <= 36'b000011001010111110001000111100111110;
		ram[565] <= 36'b000011001110110001111100111100111011;
		ram[566] <= 36'b000011010010100101100010111100110111;
		ram[567] <= 36'b000011010110011000111010111100110100;
		ram[568] <= 36'b000011011010001100000100111100110000;
		ram[569] <= 36'b000011011101111111000000111100101101;
		ram[570] <= 36'b000011100001110001110000111100101010;
		ram[571] <= 36'b000011100101100100010000111100100110;
		ram[572] <= 36'b000011101001010110100100111100100011;
		ram[573] <= 36'b000011101101001000101010111100011111;
		ram[574] <= 36'b000011110000111010100010111100011100;
		ram[575] <= 36'b000011110100101100001110111100011001;
		ram[576] <= 36'b000011111000011101101100111100010101;
		ram[577] <= 36'b000011111100001110111100111100010010;
		ram[578] <= 36'b000100000000000000000000111100001111;
		ram[579] <= 36'b000100000011110000110100111100001011;
		ram[580] <= 36'b000100000111100001011100111100001000;
		ram[581] <= 36'b000100001011010001111000111100000101;
		ram[582] <= 36'b000100001111000010000110111100000001;
		ram[583] <= 36'b000100010010110010000110111011111110;
		ram[584] <= 36'b000100010110100001111010111011111011;
		ram[585] <= 36'b000100011010010001100000111011110111;
		ram[586] <= 36'b000100011110000000111000111011110100;
		ram[587] <= 36'b000100100001110000000110111011110001;
		ram[588] <= 36'b000100100101011111000100111011101110;
		ram[589] <= 36'b000100101001001101110110111011101010;
		ram[590] <= 36'b000100101100111100011100111011100111;
		ram[591] <= 36'b000100110000101010110100111011100100;
		ram[592] <= 36'b000100110100011000111110111011100001;
		ram[593] <= 36'b000100111000000110111110111011011101;
		ram[594] <= 36'b000100111011110100101110111011011010;
		ram[595] <= 36'b000100111111100010010100111011010111;
		ram[596] <= 36'b000101000011001111101100111011010100;
		ram[597] <= 36'b000101000110111100110110111011010001;
		ram[598] <= 36'b000101001010101001110110111011001110;
		ram[599] <= 36'b000101001110010110100110111011001010;
		ram[600] <= 36'b000101010010000011001100111011000111;
		ram[601] <= 36'b000101010101101111100100111011000100;
		ram[602] <= 36'b000101011001011011110000111011000001;
		ram[603] <= 36'b000101011101000111110000111010111110;
		ram[604] <= 36'b000101100000110011100100111010111011;
		ram[605] <= 36'b000101100100011111001010111010111000;
		ram[606] <= 36'b000101101000001010100100111010110100;
		ram[607] <= 36'b000101101011110101110010111010110001;
		ram[608] <= 36'b000101101111100000110010111010101110;
		ram[609] <= 36'b000101110011001011101000111010101011;
		ram[610] <= 36'b000101110110110110010000111010101000;
		ram[611] <= 36'b000101111010100000101100111010100101;
		ram[612] <= 36'b000101111110001010111100111010100010;
		ram[613] <= 36'b000110000001110101000000111010011111;
		ram[614] <= 36'b000110000101011110110110111010011100;
		ram[615] <= 36'b000110001001001000100010111010011001;
		ram[616] <= 36'b000110001100110010000010111010010110;
		ram[617] <= 36'b000110010000011011010100111010010011;
		ram[618] <= 36'b000110010100000100011010111010010000;
		ram[619] <= 36'b000110010111101101010110111010001101;
		ram[620] <= 36'b000110011011010110000100111010001010;
		ram[621] <= 36'b000110011110111110101000111010000111;
		ram[622] <= 36'b000110100010100110111110111010000100;
		ram[623] <= 36'b000110100110001111001010111010000001;
		ram[624] <= 36'b000110101001110111001000111001111110;
		ram[625] <= 36'b000110101101011110111100111001111011;
		ram[626] <= 36'b000110110001000110100010111001111000;
		ram[627] <= 36'b000110110100101101111110111001110101;
		ram[628] <= 36'b000110111000010101001110111001110010;
		ram[629] <= 36'b000110111011111100010000111001101111;
		ram[630] <= 36'b000110111111100011001000111001101100;
		ram[631] <= 36'b000111000011001001110110111001101001;
		ram[632] <= 36'b000111000110110000010110111001100110;
		ram[633] <= 36'b000111001010010110101010111001100011;
		ram[634] <= 36'b000111001101111100110100111001100000;
		ram[635] <= 36'b000111010001100010110010111001011101;
		ram[636] <= 36'b000111010101001000100100111001011011;
		ram[637] <= 36'b000111011000101110001010111001011000;
		ram[638] <= 36'b000111011100010011100110111001010101;
		ram[639] <= 36'b000111011111111000110100111001010010;
		ram[640] <= 36'b000111100011011101111000111001001111;
		ram[641] <= 36'b000111100111000010110010111001001100;
		ram[642] <= 36'b000111101010100111011110111001001001;
		ram[643] <= 36'b000111101110001100000000111001000111;
		ram[644] <= 36'b000111110001110000010110111001000100;
		ram[645] <= 36'b000111110101010100100010111001000001;
		ram[646] <= 36'b000111111000111000100010111000111110;
		ram[647] <= 36'b000111111100011100010110111000111011;
		ram[648] <= 36'b001000000000000000000000111000111000;
		ram[649] <= 36'b001000000011100011011100111000110110;
		ram[650] <= 36'b001000000111000110110000111000110011;
		ram[651] <= 36'b001000001010101001111000111000110000;
		ram[652] <= 36'b001000001110001100110100111000101101;
		ram[653] <= 36'b001000010001101111100100111000101010;
		ram[654] <= 36'b001000010101010010001010111000101000;
		ram[655] <= 36'b001000011000110100100110111000100101;
		ram[656] <= 36'b001000011100010110110110111000100010;
		ram[657] <= 36'b001000011111111000111100111000011111;
		ram[658] <= 36'b001000100011011010110100111000011101;
		ram[659] <= 36'b001000100110111100100100111000011010;
		ram[660] <= 36'b001000101010011110001000111000010111;
		ram[661] <= 36'b001000101101111111100010111000010100;
		ram[662] <= 36'b001000110001100000110000111000010010;
		ram[663] <= 36'b001000110101000001110010111000001111;
		ram[664] <= 36'b001000111000100010101100111000001100;
		ram[665] <= 36'b001000111100000011011000111000001010;
		ram[666] <= 36'b001000111111100011111100111000000111;
		ram[667] <= 36'b001001000011000100010100111000000100;
		ram[668] <= 36'b001001000110100100100000111000000001;
		ram[669] <= 36'b001001001010000100100100110111111111;
		ram[670] <= 36'b001001001101100100011010110111111100;
		ram[671] <= 36'b001001010001000100001000110111111001;
		ram[672] <= 36'b001001010100100011101010110111110111;
		ram[673] <= 36'b001001011000000011000010110111110100;
		ram[674] <= 36'b001001011011100010010000110111110001;
		ram[675] <= 36'b001001011111000001010010110111101111;
		ram[676] <= 36'b001001100010100000001010110111101100;
		ram[677] <= 36'b001001100101111110111000110111101010;
		ram[678] <= 36'b001001101001011101011010110111100111;
		ram[679] <= 36'b001001101100111011110100110111100100;
		ram[680] <= 36'b001001110000011010000010110111100010;
		ram[681] <= 36'b001001110011111000000100110111011111;
		ram[682] <= 36'b001001110111010101111110110111011100;
		ram[683] <= 36'b001001111010110011101100110111011010;
		ram[684] <= 36'b001001111110010001010000110111010111;
		ram[685] <= 36'b001010000001101110101010110111010101;
		ram[686] <= 36'b001010000101001011111010110111010010;
		ram[687] <= 36'b001010001000101001000000110111010000;
		ram[688] <= 36'b001010001100000101111010110111001101;
		ram[689] <= 36'b001010001111100010101100110111001010;
		ram[690] <= 36'b001010010010111111010010110111001000;
		ram[691] <= 36'b001010010110011011101110110111000101;
		ram[692] <= 36'b001010011001111000000000110111000011;
		ram[693] <= 36'b001010011101010100001000110111000000;
		ram[694] <= 36'b001010100000110000000110110110111110;
		ram[695] <= 36'b001010100100001011111010110110111011;
		ram[696] <= 36'b001010100111100111100010110110111001;
		ram[697] <= 36'b001010101011000011000010110110110110;
		ram[698] <= 36'b001010101110011110011000110110110100;
		ram[699] <= 36'b001010110001111001100010110110110001;
		ram[700] <= 36'b001010110101010100100100110110101111;
		ram[701] <= 36'b001010111000101111011010110110101100;
		ram[702] <= 36'b001010111100001010001000110110101010;
		ram[703] <= 36'b001010111111100100101100110110100111;
		ram[704] <= 36'b001011000010111111000100110110100101;
		ram[705] <= 36'b001011000110011001010100110110100010;
		ram[706] <= 36'b001011001001110011011010110110100000;
		ram[707] <= 36'b001011001101001101010100110110011101;
		ram[708] <= 36'b001011010000100111000110110110011011;
		ram[709] <= 36'b001011010100000000101110110110011000;
		ram[710] <= 36'b001011010111011010001100110110010110;
		ram[711] <= 36'b001011011010110011100000110110010011;
		ram[712] <= 36'b001011011110001100101100110110010001;
		ram[713] <= 36'b001011100001100101101100110110001110;
		ram[714] <= 36'b001011100100111110100100110110001100;
		ram[715] <= 36'b001011101000010111010000110110001010;
		ram[716] <= 36'b001011101011101111110100110110000111;
		ram[717] <= 36'b001011101111001000001110110110000101;
		ram[718] <= 36'b001011110010100000011110110110000010;
		ram[719] <= 36'b001011110101111000100100110110000000;
		ram[720] <= 36'b001011111001010000100010110101111110;
		ram[721] <= 36'b001011111100101000010110110101111011;
		ram[722] <= 36'b001100000000000000000000110101111001;
		ram[723] <= 36'b001100000011010111100000110101110110;
		ram[724] <= 36'b001100000110101110110110110101110100;
		ram[725] <= 36'b001100001010000110000100110101110010;
		ram[726] <= 36'b001100001101011101000110110101101111;
		ram[727] <= 36'b001100010000110100000010110101101101;
		ram[728] <= 36'b001100010100001010110010110101101011;
		ram[729] <= 36'b001100010111100001011010110101101000;
		ram[730] <= 36'b001100011010110111111000110101100110;
		ram[731] <= 36'b001100011110001110001100110101100011;
		ram[732] <= 36'b001100100001100100011000110101100001;
		ram[733] <= 36'b001100100100111010011000110101011111;
		ram[734] <= 36'b001100101000010000010010110101011100;
		ram[735] <= 36'b001100101011100110000000110101011010;
		ram[736] <= 36'b001100101110111011100110110101011000;
		ram[737] <= 36'b001100110010010001000010110101010101;
		ram[738] <= 36'b001100110101100110010110110101010011;
		ram[739] <= 36'b001100111000111011100000110101010001;
		ram[740] <= 36'b001100111100010000100010110101001111;
		ram[741] <= 36'b001100111111100101011000110101001100;
		ram[742] <= 36'b001101000010111010001000110101001010;
		ram[743] <= 36'b001101000110001110101100110101001000;
		ram[744] <= 36'b001101001001100011001000110101000101;
		ram[745] <= 36'b001101001100110111011100110101000011;
		ram[746] <= 36'b001101010000001011100110110101000001;
		ram[747] <= 36'b001101010011011111100110110100111111;
		ram[748] <= 36'b001101010110110011011110110100111100;
		ram[749] <= 36'b001101011010000111001100110100111010;
		ram[750] <= 36'b001101011101011010110010110100111000;
		ram[751] <= 36'b001101100000101110001110110100110110;
		ram[752] <= 36'b001101100100000001100010110100110011;
		ram[753] <= 36'b001101100111010100101100110100110001;
		ram[754] <= 36'b001101101010100111101110110100101111;
		ram[755] <= 36'b001101101101111010100110110100101101;
		ram[756] <= 36'b001101110001001101010110110100101010;
		ram[757] <= 36'b001101110100011111111110110100101000;
		ram[758] <= 36'b001101110111110010011100110100100110;
		ram[759] <= 36'b001101111011000100110000110100100100;
		ram[760] <= 36'b001101111110010110111100110100100001;
		ram[761] <= 36'b001110000001101001000000110100011111;
		ram[762] <= 36'b001110000100111010111010110100011101;
		ram[763] <= 36'b001110001000001100101100110100011011;
		ram[764] <= 36'b001110001011011110010100110100011001;
		ram[765] <= 36'b001110001110101111110100110100010110;
		ram[766] <= 36'b001110010010000001001100110100010100;
		ram[767] <= 36'b001110010101010010011010110100010010;
		ram[768] <= 36'b001110011000100011100000110100010000;
		ram[769] <= 36'b001110011011110100011110110100001110;
		ram[770] <= 36'b001110011111000101010010110100001100;
		ram[771] <= 36'b001110100010010101111110110100001001;
		ram[772] <= 36'b001110100101100110100000110100000111;
		ram[773] <= 36'b001110101000110110111100110100000101;
		ram[774] <= 36'b001110101100000111001100110100000011;
		ram[775] <= 36'b001110101111010111010110110100000001;
		ram[776] <= 36'b001110110010100111010110110011111111;
		ram[777] <= 36'b001110110101110111001110110011111100;
		ram[778] <= 36'b001110111001000110111110110011111010;
		ram[779] <= 36'b001110111100010110100110110011111000;
		ram[780] <= 36'b001110111111100110000100110011110110;
		ram[781] <= 36'b001111000010110101011010110011110100;
		ram[782] <= 36'b001111000110000100101000110011110010;
		ram[783] <= 36'b001111001001010011101100110011110000;
		ram[784] <= 36'b001111001100100010101000110011101110;
		ram[785] <= 36'b001111001111110001011100110011101011;
		ram[786] <= 36'b001111010011000000001000110011101001;
		ram[787] <= 36'b001111010110001110101100110011100111;
		ram[788] <= 36'b001111011001011101000110110011100101;
		ram[789] <= 36'b001111011100101011011000110011100011;
		ram[790] <= 36'b001111011111111001100010110011100001;
		ram[791] <= 36'b001111100011000111100100110011011111;
		ram[792] <= 36'b001111100110010101011110110011011101;
		ram[793] <= 36'b001111101001100011010000110011011011;
		ram[794] <= 36'b001111101100110000111000110011011001;
		ram[795] <= 36'b001111101111111110011000110011010111;
		ram[796] <= 36'b001111110011001011110000110011010101;
		ram[797] <= 36'b001111110110011001000000110011010010;
		ram[798] <= 36'b001111111001100110001000110011010000;
		ram[799] <= 36'b001111111100110011001000110011001110;
		ram[800] <= 36'b010000000000000000000000110011001100;
		ram[801] <= 36'b010000000011001100101110110011001010;
		ram[802] <= 36'b010000000110011001010110110011001000;
		ram[803] <= 36'b010000001001100101110100110011000110;
		ram[804] <= 36'b010000001100110010001010110011000100;
		ram[805] <= 36'b010000001111111110011000110011000010;
		ram[806] <= 36'b010000010011001010100000110011000000;
		ram[807] <= 36'b010000010110010110011110110010111110;
		ram[808] <= 36'b010000011001100010010100110010111100;
		ram[809] <= 36'b010000011100101110000010110010111010;
		ram[810] <= 36'b010000011111111001101000110010111000;
		ram[811] <= 36'b010000100011000101000110110010110110;
		ram[812] <= 36'b010000100110010000011100110010110100;
		ram[813] <= 36'b010000101001011011101010110010110010;
		ram[814] <= 36'b010000101100100110110000110010110000;
		ram[815] <= 36'b010000101111110001101110110010101110;
		ram[816] <= 36'b010000110010111100100100110010101100;
		ram[817] <= 36'b010000110110000111010010110010101010;
		ram[818] <= 36'b010000111001010001111000110010101000;
		ram[819] <= 36'b010000111100011100010110110010100110;
		ram[820] <= 36'b010000111111100110101100110010100100;
		ram[821] <= 36'b010001000010110000111100110010100010;
		ram[822] <= 36'b010001000101111011000010110010100000;
		ram[823] <= 36'b010001001001000101000000110010011110;
		ram[824] <= 36'b010001001100001110111000110010011100;
		ram[825] <= 36'b010001001111011000100110110010011010;
		ram[826] <= 36'b010001010010100010001110110010011000;
		ram[827] <= 36'b010001010101101011101100110010010110;
		ram[828] <= 36'b010001011000110101000100110010010100;
		ram[829] <= 36'b010001011011111110010100110010010010;
		ram[830] <= 36'b010001011111000111011100110010010001;
		ram[831] <= 36'b010001100010010000011100110010001111;
		ram[832] <= 36'b010001100101011001010100110010001101;
		ram[833] <= 36'b010001101000100010000110110010001011;
		ram[834] <= 36'b010001101011101010101110110010001001;
		ram[835] <= 36'b010001101110110011010000110010000111;
		ram[836] <= 36'b010001110001111011101010110010000101;
		ram[837] <= 36'b010001110101000011111100110010000011;
		ram[838] <= 36'b010001111000001100000110110010000001;
		ram[839] <= 36'b010001111011010100001010110001111111;
		ram[840] <= 36'b010001111110011100000100110001111101;
		ram[841] <= 36'b010010000001100011111000110001111011;
		ram[842] <= 36'b010010000100101011100100110001111010;
		ram[843] <= 36'b010010000111110011001000110001111000;
		ram[844] <= 36'b010010001010111010100100110001110110;
		ram[845] <= 36'b010010001110000001111010110001110100;
		ram[846] <= 36'b010010010001001001001000110001110010;
		ram[847] <= 36'b010010010100010000001110110001110000;
		ram[848] <= 36'b010010010111010111001100110001101110;
		ram[849] <= 36'b010010011010011110000100110001101100;
		ram[850] <= 36'b010010011101100100110100110001101010;
		ram[851] <= 36'b010010100000101011011100110001101001;
		ram[852] <= 36'b010010100011110001111100110001100111;
		ram[853] <= 36'b010010100110111000010100110001100101;
		ram[854] <= 36'b010010101001111110100110110001100011;
		ram[855] <= 36'b010010101101000100110010110001100001;
		ram[856] <= 36'b010010110000001010110100110001011111;
		ram[857] <= 36'b010010110011010000110000110001011101;
		ram[858] <= 36'b010010110110010110100100110001011100;
		ram[859] <= 36'b010010111001011100010000110001011010;
		ram[860] <= 36'b010010111100100001110110110001011000;
		ram[861] <= 36'b010010111111100111010100110001010110;
		ram[862] <= 36'b010011000010101100101010110001010100;
		ram[863] <= 36'b010011000101110001111010110001010010;
		ram[864] <= 36'b010011001000110111000010110001010001;
		ram[865] <= 36'b010011001011111100000010110001001111;
		ram[866] <= 36'b010011001111000000111100110001001101;
		ram[867] <= 36'b010011010010000101101110110001001011;
		ram[868] <= 36'b010011010101001010011010110001001001;
		ram[869] <= 36'b010011011000001110111100110001001000;
		ram[870] <= 36'b010011011011010011011010110001000110;
		ram[871] <= 36'b010011011110010111101110110001000100;
		ram[872] <= 36'b010011100001011011111100110001000010;
		ram[873] <= 36'b010011100100100000000100110001000000;
		ram[874] <= 36'b010011100111100100000100110000111111;
		ram[875] <= 36'b010011101010100111111100110000111101;
		ram[876] <= 36'b010011101101101011101100110000111011;
		ram[877] <= 36'b010011110000101111011000110000111001;
		ram[878] <= 36'b010011110011110010111010110000110111;
		ram[879] <= 36'b010011110110110110010110110000110110;
		ram[880] <= 36'b010011111001111001101010110000110100;
		ram[881] <= 36'b010011111100111100111000110000110010;
		ram[882] <= 36'b010100000000000000000000110000110000;
		ram[883] <= 36'b010100000011000010111110110000101110;
		ram[884] <= 36'b010100000110000101110110110000101101;
		ram[885] <= 36'b010100001001001000101000110000101011;
		ram[886] <= 36'b010100001100001011010010110000101001;
		ram[887] <= 36'b010100001111001101110110110000100111;
		ram[888] <= 36'b010100010010010000010010110000100110;
		ram[889] <= 36'b010100010101010010101000110000100100;
		ram[890] <= 36'b010100011000010100110110110000100010;
		ram[891] <= 36'b010100011011010110111110110000100000;
		ram[892] <= 36'b010100011110011000111110110000011111;
		ram[893] <= 36'b010100100001011010111000110000011101;
		ram[894] <= 36'b010100100100011100101010110000011011;
		ram[895] <= 36'b010100100111011110010110110000011010;
		ram[896] <= 36'b010100101010011111111010110000011000;
		ram[897] <= 36'b010100101101100001011000110000010110;
		ram[898] <= 36'b010100110000100010101110110000010100;
		ram[899] <= 36'b010100110011100011111110110000010011;
		ram[900] <= 36'b010100110110100101001000110000010001;
		ram[901] <= 36'b010100111001100110001010110000001111;
		ram[902] <= 36'b010100111100100111000100110000001101;
		ram[903] <= 36'b010100111111100111111000110000001100;
		ram[904] <= 36'b010101000010101000100110110000001010;
		ram[905] <= 36'b010101000101101001001110110000001000;
		ram[906] <= 36'b010101001000101001101110110000000111;
		ram[907] <= 36'b010101001011101010000110110000000101;
		ram[908] <= 36'b010101001110101010011000110000000011;
		ram[909] <= 36'b010101010001101010100100110000000010;
		ram[910] <= 36'b010101010100101010101010110000000000;
		ram[911] <= 36'b010101010111101010101000101111111110;
		ram[912] <= 36'b010101011010101010100000101111111101;
		ram[913] <= 36'b010101011101101010010000101111111011;
		ram[914] <= 36'b010101100000101001111010101111111001;
		ram[915] <= 36'b010101100011101001011100101111110111;
		ram[916] <= 36'b010101100110101000111010101111110110;
		ram[917] <= 36'b010101101001101000010000101111110100;
		ram[918] <= 36'b010101101100100111011110101111110010;
		ram[919] <= 36'b010101101111100110100110101111110001;
		ram[920] <= 36'b010101110010100101101000101111101111;
		ram[921] <= 36'b010101110101100100100100101111101101;
		ram[922] <= 36'b010101111000100011011000101111101100;
		ram[923] <= 36'b010101111011100010000110101111101010;
		ram[924] <= 36'b010101111110100000101110101111101001;
		ram[925] <= 36'b010110000001011111001110101111100111;
		ram[926] <= 36'b010110000100011101101000101111100101;
		ram[927] <= 36'b010110000111011011111100101111100100;
		ram[928] <= 36'b010110001010011010001010101111100010;
		ram[929] <= 36'b010110001101011000010000101111100000;
		ram[930] <= 36'b010110010000010110010000101111011111;
		ram[931] <= 36'b010110010011010100001010101111011101;
		ram[932] <= 36'b010110010110010001111100101111011011;
		ram[933] <= 36'b010110011001001111101000101111011010;
		ram[934] <= 36'b010110011100001101001110101111011000;
		ram[935] <= 36'b010110011111001010101110101111010111;
		ram[936] <= 36'b010110100010001000000110101111010101;
		ram[937] <= 36'b010110100101000101011000101111010011;
		ram[938] <= 36'b010110101000000010100100101111010010;
		ram[939] <= 36'b010110101010111111101010101111010000;
		ram[940] <= 36'b010110101101111100101000101111001110;
		ram[941] <= 36'b010110110000111001100010101111001101;
		ram[942] <= 36'b010110110011110110010100101111001011;
		ram[943] <= 36'b010110110110110011000000101111001010;
		ram[944] <= 36'b010110111001101111100100101111001000;
		ram[945] <= 36'b010110111100101100000100101111000110;
		ram[946] <= 36'b010110111111101000011100101111000101;
		ram[947] <= 36'b010111000010100100101110101111000011;
		ram[948] <= 36'b010111000101100000111010101111000010;
		ram[949] <= 36'b010111001000011101000000101111000000;
		ram[950] <= 36'b010111001011011001000000101110111110;
		ram[951] <= 36'b010111001110010100111000101110111101;
		ram[952] <= 36'b010111010001010000101010101110111011;
		ram[953] <= 36'b010111010100001100010110101110111010;
		ram[954] <= 36'b010111010111000111111100101110111000;
		ram[955] <= 36'b010111011010000011011100101110110111;
		ram[956] <= 36'b010111011100111110110110101110110101;
		ram[957] <= 36'b010111011111111010001000101110110011;
		ram[958] <= 36'b010111100010110101010110101110110010;
		ram[959] <= 36'b010111100101110000011100101110110000;
		ram[960] <= 36'b010111101000101011011100101110101111;
		ram[961] <= 36'b010111101011100110010110101110101101;
		ram[962] <= 36'b010111101110100001001010101110101100;
		ram[963] <= 36'b010111110001011011111000101110101010;
		ram[964] <= 36'b010111110100010110100000101110101001;
		ram[965] <= 36'b010111110111010001000000101110100111;
		ram[966] <= 36'b010111111010001011011100101110100101;
		ram[967] <= 36'b010111111101000101110000101110100100;
		ram[968] <= 36'b011000000000000000000000101110100010;
		ram[969] <= 36'b011000000010111010001000101110100001;
		ram[970] <= 36'b011000000101110100001010101110011111;
		ram[971] <= 36'b011000001000101110000110101110011110;
		ram[972] <= 36'b011000001011100111111100101110011100;
		ram[973] <= 36'b011000001110100001101100101110011011;
		ram[974] <= 36'b011000010001011011010110101110011001;
		ram[975] <= 36'b011000010100010100111010101110011000;
		ram[976] <= 36'b011000010111001110011000101110010110;
		ram[977] <= 36'b011000011010000111110000101110010101;
		ram[978] <= 36'b011000011101000001000010101110010011;
		ram[979] <= 36'b011000011111111010001100101110010010;
		ram[980] <= 36'b011000100010110011010010101110010000;
		ram[981] <= 36'b011000100101101100010010101110001111;
		ram[982] <= 36'b011000101000100101001100101110001101;
		ram[983] <= 36'b011000101011011101111110101110001100;
		ram[984] <= 36'b011000101110010110101100101110001010;
		ram[985] <= 36'b011000110001001111010100101110001001;
		ram[986] <= 36'b011000110100000111110100101110000111;
		ram[987] <= 36'b011000110111000000010000101110000110;
		ram[988] <= 36'b011000111001111000100110101110000100;
		ram[989] <= 36'b011000111100110000110100101110000011;
		ram[990] <= 36'b011000111111101000111110101110000001;
		ram[991] <= 36'b011001000010100001000010101110000000;
		ram[992] <= 36'b011001000101011001000000101101111110;
		ram[993] <= 36'b011001001000010000110110101101111101;
		ram[994] <= 36'b011001001011001000101000101101111011;
		ram[995] <= 36'b011001001110000000010100101101111010;
		ram[996] <= 36'b011001010000110111111010101101111000;
		ram[997] <= 36'b011001010011101111011010101101110111;
		ram[998] <= 36'b011001010110100110110100101101110101;
		ram[999] <= 36'b011001011001011110001000101101110100;
		ram[1000] <= 36'b011001011100010101011000101101110010;
		ram[1001] <= 36'b011001011111001100100000101101110001;
		ram[1002] <= 36'b011001100010000011100010101101101111;
		ram[1003] <= 36'b011001100100111010100000101101101110;
		ram[1004] <= 36'b011001100111110001010110101101101101;
		ram[1005] <= 36'b011001101010101000001000101101101011;
		ram[1006] <= 36'b011001101101011110110010101101101010;
		ram[1007] <= 36'b011001110000010101011000101101101000;
		ram[1008] <= 36'b011001110011001011111000101101100111;
		ram[1009] <= 36'b011001110110000010010010101101100101;
		ram[1010] <= 36'b011001111000111000100110101101100100;
		ram[1011] <= 36'b011001111011101110110100101101100010;
		ram[1012] <= 36'b011001111110100100111100101101100001;
		ram[1013] <= 36'b011010000001011011000000101101011111;
		ram[1014] <= 36'b011010000100010000111100101101011110;
		ram[1015] <= 36'b011010000111000110110100101101011101;
		ram[1016] <= 36'b011010001001111100100110101101011011;
		ram[1017] <= 36'b011010001100110010010010101101011010;
		ram[1018] <= 36'b011010001111100111111000101101011000;
		ram[1019] <= 36'b011010010010011101011000101101010111;
		ram[1020] <= 36'b011010010101010010110100101101010101;
		ram[1021] <= 36'b011010011000001000001000101101010100;
		ram[1022] <= 36'b011010011010111101011000101101010011;
		ram[1023] <= 36'b011010011101110010100010101101010001;
    end
    ram_read <= ram[op[23:14]];
    exp2 <= op[30:23] >> 1'b1;
    res <= op[13:0];
end

always @(posedge clk) begin
    grad_mul_res <= ram_grad * res;
    exp3 <= exp2;
    frac <= ram_main;
end

wire [23:0] grad_mul_res_need;
assign grad_mul_res_need = {1'b0, grad_mul_res[26:4]};
wire [23:0] result_1;//[23]は必ず1になるはず：デバッグ用
assign result_1 = frac + grad_mul_res_need;

wire [23:0] result_plus1_1;
assign result_plus1_1 = result_1 + 24'd1;

always @(posedge clk) begin
    if (ready) begin
        ready <= 1'b0;
    end
    if (grad_mul_res[3]) begin//精度が大丈夫そうなら消したほうが早いかも
        result <= {1'b0, exp3, result_plus1_1[22:0]};
        ready <= 1'b1;
    end else begin
        result <= {1'b0, exp3, result_1[22:0]};
        ready <= 1'b1;
    end
end
endmodule
`default_nettype wire